��[ M a i n ]  
 C a p t i o n 	 = " I n s t a l l   N a v i   [ % P R O D U C T _ N A M E % ] "  
 B T N _ N e x t 	 = " N � s t a "  
 B T N _ B a c k 	 = " B a k � t "  
 B T N _ I n s t a l l 	 = " I n s t a l l e r a "  
 B T N _ C a n c e l 	 = " A v b r y t "  
 B T N _ F i n i s h 	 = " S l u t f � r "  
 B T N _ S k i p 	 = " H o p p a   � v e r "  
 B T N _ A p p l y 	 = " V e r k s t � l l "  
 B T N _ R e g i s t 	 = " R e g i s t r e r a "  
 B T N _ R e s t a r t 	 = " M o d e l l � t e r s t � l l n i n g "  
 P D M _ L a n g u a g e 	 = " S p r � k "  
 D L G _ C a n c e l 	 = " � r   d u   s � k e r   p �   a t t   d u   v i l l   a v b r y t a ? "  
 L B L _ P r i n t e r 	 = " S k r i v a r e "  
 L B L _ S c a n n e r 	 = " S k a n n e r "  
 L B L _ W i f i 	 = " W i - F i - a n s l u t n i n g "  
 L B L _ R e c o m m e n d e d 	 = " ( R e k o m m e n d e r a s ) "  
  
 [ S t a r t M e n u ]  
 T I T L E 	 = " I n s t a l l   N a v i "  
 S U B _ T i t l e 	 = " "  
 L N K _ S t a r t 	 = " S t a r t   o c h   a n s l u t n i n g "  
 H L P _ S t a r t 	 = " K l i c k a   h � r   n � r   d u   v i l l   s t a r t a   i n s t a l l a t i o n s p r o c e s s e n ,   i n s t a l l e r a   p r o g r a m v a r a n   o c h   k o n f i g u r e r a   n � t v e r k s i n s t � l l n i n g a r . "  
 L N K _ G u i d e 	 = " E n d a s t   f � r   s y s t e m a d m i n i s t r a t � r e r "  
 H L P _ G u i d e 	 = " K l i c k a   h � r   o m   d u   v i l l   v i s a   s k r i v a r e n s   h a n d b o k   o m   m a s k i n v a r u i n s t a l l a t i o n   ( P D F )   o c h   a n d r a   a d m i n i s t r a t i v a   i n s t � l l n i n g a r . "  
 L N K _ M o d e l 	 = " V � l j   d i n   p r o d u k t "  
 H L P _ M o d e l 	 = " M a r k e r a   p r o d u k t e n   i   l i s t a n . "  
 L N K _ M a n u a l 	 = " I n f o r m a t i o n   f � r   h a n d b � c k e r   o c h   p r o g r a m "  
 H L P _ M a n u a l 	 = " K l i c k a   h � r   f � r   a t t   f �   i n f o r m a t i o n   o m   h a n d b � c k e r ,   d e   v a n l i g a s t e   p r o g r a m m e n   s � s o m   s k r i v a r d r i v r u t i n e r   o c h   s � k v � g a r   t i l l   d e s s a   p r o g r a m   s o m   f i n n s   p �   p r o g r a m v a r a n s   c d - s k i v a   s �   a t t   d u   k a n   i n s t a l l e r a   d e m   m a n u e l l t . "  
  
 [ S e l e c t M o d e l ]  
 T I T L E = " V � l j   d i n   p r o d u k t "  
 T X T _ B o d y = " M a r k e r a   p r o d u k t e n   i   l i s t a n . "  
  
 [ F o r A d m i n ]  
 T I T L E 	 = " E n d a s t   f � r   s y s t e m a d m i n i s t r a t � r e r "  
 S U B _ T i t l e 	 = " "  
 B T N _ H S G 	 = " H a n d b o k   f � r   m a s k i n v a r u i n s t a l l a t i o n "  
  
 [ V i e w M a n u a l ]  
 T I T L E 	 = " I n f o r m a t i o n   f � r   h a n d b � c k e r   o c h   p r o g r a m "  
 S U B _ T i t l e 	 = " "  
 B T N _ F o l d e r 	 = " H a n d b � c k e r "  
  
 [ L i c e n s e A a g r e e m e n t ]  
 T I T L E 	 = " L i c e n s a v t a l "  
 S U B _ T i t l e 	 = " L � s   l i c e n s a v t a l e t   n o g a . "  
 L N K _ O p t i o n 	 = " A l t e r n a t i v   f � r   i n s t a l l a t i o n   a v   p r o g r a m v a r a "  
 C B X _ A g r e e 	 = " J a g   g o d k � n n e r   l i c e n s a v t a l e t . "  
 I T M _ L a n g u a g e 	 = " S p r � k "  
  
 [ S y s t e m C h e c k ]  
 T I T L E 	 = " F � r b e r e d e r   i n s t a l l a t i o n "  
 S U B _ T i t l e 	 = " "  
 T X T _ C h e c k P C 	 = " F � r b e r e d e r   i n s t a l l a t i o n   . . .   v � n t a . "  
 T X T _ C h e c k N W 	 = " F � r b e r e d e r   i n s t a l l a t i o n   . . .   v � n t a . "  
  
 [ S e l e c t D r i v e r M e n u ]  
 T I T L E 	 = " V � l j   s k r i v a r d r i v r u t i n "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " V � l j   e n   s k r i v a r d r i v r u t i n   s o m   d u   v i l l   i n s t a l l e r a . "  
 R B T _ G D I 	 = " S k r i v a r d r i v r u t i n e n   G D I   ( G r a p h i c s   D e v i c e   I n t e r f a c e ) "  
 H L P _ G D I 	 = " M e d   s k r i v a r d r i v r u t i n e n   k o m m e r   p r o g r a m v a r a n   s o m   m a x i m e r a r   s k r i v a r e n s   f u n k t i o n   o c h   k o n f i g u r e r a r   n � t v e r k s i n s t � l l n i n g a r   o c k s �   a t t   i n s t a l l e r a s . "  
 R B T _ A D D 	 = " A n d r a   s k r i v a r d r i v r u t i n e r   � n   o v a n . "  
 H L P _ A D D 	 = " K l i c k a   h � r   o m   d u   b a r a   v i l l   i n s t a l l e r a   P C L - s k r i v a r d r i v r u t i n e n   e l l e r   P S 3 - s k r i v a r d r i v r u t i n e n . "  
  
 [ D o w n l o a d E a c h D r i v e r ]  
 T I T L E 	 = " H � m t a   d r i v r u t i n e r   o c h   p r o g r a m "  
 T X T _ B o d y 	 = " V � l j   s k r i v a r d r i v r u t i n e n   e l l e r   p r o g r a m v a r a n   s o m   d u   v i l l   h � m t a . "  
 L N K _ P C L 	 = " P C L - s k r i v a r d r i v r u t i n e n "  
 L N K _ P S 3 	 = " P S 3   ( P o s t S c r i p t 3 ) - s k r i v a r d r i v r u t i n e n "  
 L N K _ E N C 	 = " E p s o n N e t   C o n f i g "  
 C A U T I O N 	 = " V i s s a   f u n k t i o n e r   � r   i n t e   t i l l g � n g l i g a   m e d   d e s s a   d r i v r u t i n e r .   O m   d u   v i l l   a n v � n d a   a l l a   s k r i v a r e n s   f u n k t i o n e r ,   g �   t i l l b a k a   t i l l   f � r e g � e n d e   s k � r m   o c h   i n s t a l l e r a   G D I - s k r i v a r d r i v r u t i n e n . "  
  
 [ I n s t a l l O p t i o n ]  
 T I T L E 	 = " A l t e r n a t i v   f � r   i n s t a l l a t i o n   a v   p r o g r a m v a r a "  
 S U B _ T i t l e 	 = " V � l j   v i l k a   i n s t a l l a t i o n s a l t e r n a t i v   d u   v i l l   a n v � n d a . "  
 T X T _ B o d y 	 = " "  
 C B X _ L a t e s t 	 = " I n s t a l l e r a   d e n   s e n a s t e   v e r s i o n e n   % R E C O M M E N D E D % "  
 H L P _ L a t e s t 	 = " I n s t a l l e r a   d e n   s e n a s t e   v e r s i o n e n   a v   d r i v r u t i n e n   f r � n   E p s o n s   w e b b p l a t s . "  
 C B X _ S t a t u s 	 = " � v e r v a k n i n g   a v   p r o d u k t s t a t u s   o c h   a u t o m a t i s k a   u p p d a t e r i n g a r   % R E C O M M E N D E D % "  
 H L P _ S t a t u s 	 = " A n v � n d s   f � r   a t t   a u t o m a t i s k t   k o n t r o l l e r a   o c h   i n s t a l l e r a   d e   s e n a s t e   u p p d a t e r i n g a r n a   f � r   p r o d u k t e n .   I n g a   p e r s o n u p p g i f t e r   k o m m e r   a t t   h � m t a s . "  
  
 [ R e I n s t a l l ]  
 T I T L E 	 = " V � l j   p r o g r a m v a r u i n s t a l l a t i o n "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " I n s t a l l a t i o n s p r o g r a m m e t   h a r   u p p t � c k t   a t t   % P R O D U C T % n   r e d a n   h a r   i n s t a l l e r a t s   p �   d a t o r n . \ r \ n V � l j   m e l l a n   f � l j a n d e   a l t e r n a t i v : "  
 R B T _ E s s e n t i l a l 	 = " O m i n s t a l l e r a   p r o g r a m v a r a n "  
 H L P _ E s s e n t i l a l 	 = " V � l j   d e t t a   o m   d u   v i l l   o m i n s t a l l e r a   p r o g r a m v a r a n   o c h   � n d r a   a n s l u t n i n g s i n s t � l l n i n g a r n a   f � r   % P R O D U C T % n . "  
 R B T _ A d d S o f t 	 = " I n s t a l l e r a   t i l l � m p n i n g s p r o g r a m "  
 H L P _ A d d S o f t 	 = " I n s t a l l e r a   � v r i g a   E p s o n - p r o g r a m . "  
  
 [ P r i n t e r L i s t ]  
 T I T L E 	 = " F � r s t a   i n s t a l l a t i o n e n ? "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " � r   d e t   f � r s t a   g � n g e n   d u   i n s t a l l e r a r   % P R O D U C T % n ? "  
 R B T _ F i r s t 	 = " J a ,   d e t   � r   f � r s t a   g � n g e n "  
 H L P _ F i r s t 	 = " D u   k o m m e r   b l i   g u i d a d   g e n o m   i n s t a l l a t i o n s p r o c e s s e n   f � r   % P R O D U C T % n . "  
 R B T _ A d d i n g 	 = " % P R O D U C T %   a n v � n d s   r e d a n   -   t i l l � t   d a t o r n   a t t   s k r i v a   u t "  
 H L P _ A d d i n g 	 = " V � l j   % P R O D U C T % n   f r � n   l i s t a n   n e d a n .   O m   d e n   i n t e   f i n n s   m e d   i   l i s t a n   k o n t r o l l e r a r   d u   a t t   % P R O D U C T % n   � r   p �   o c h   a n s l u t e n   t i l l   d i t t   n � t v e r k . "  
 L S T _ M o d e l 	 = " p r o d u k t "  
 L S T _ M a c A d d r e s s 	 = " M A C - a d r e s s "  
 L S T _ I P A d d r e s s 	 = " I P - a d r e s s "  
 L N K _ I P _ M A N U A L 	 = " A v a n c e r a d   k o n f i g u r a t i o n "  
  
 [ I P M a n u a l S e t u p ]  
 T I T L E 	 = " V � l j a   I P - a d r e s s   m a n u e l l t "  
 S U B _ T I T L E 	 = " "  
 T X T _ B o d y 	 = " A n g e   I P - a d r e s s   i   r u t a n   n e d a n .   % P R O D U C T % p o r t e n   k o n f i g u r e r a s   m e d   d e n   I P - a d r e s s e n . "  
 I T M _ I P 	 = " I P - a d r e s s : "  
  
 [ H a r d w a r e S e t u p ]  
 T I T L E 	 = " I n s t a l l e r a "  
 S U B _ T i t l e 	 = " "  
  
 [ I n s t a l l E s s e n t i a l ]  
 T I T L E 	 = " I n s t a l l e r a r   p r o g r a m v a r a "  
 T I T L E _ D L 	 = " N e r l a d d n i n g   E s s e n t i a l - p r o g r a m v a r a "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y _ D L 	 = " H � m t a r   . . .   % s "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   . . .   % s "  
  
 [ S e l e c t C o n n e c t ]  
 T I T L E 	 = " A n s l u t   % P R O D U C T % "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " V � l j   h u r   d u   v i l l   a n s l u t a   % P R O D U C T % n   t i l l   d a t o r n   e l l e r   t i l l   e n   a n n a n   e n h e t . "  
 R B T _ W i f i 	 = " % W I F I % "  
 R B T _ W A C 	 = " % W I F I %   % R E C O M M E N D E D % "  
 H L P _ W i f i 	 = " U p p r � t t a r   e n   t r � d l � s   a n s l u t n i n g   t i l l   % P R O D U C T % n . "  
 R B T _ L A N 	 = " E t h e r n e t - a n s l u t n i n g "  
 H L P _ L A N 	 = " V � l j   d e n n a   o m   d u   a n v � n d e r   e t t   k a b e l a n s l u t e t   n � t v e r k   o c h   v i l l   a n s l u t a   m e d   h j � l p   a v   e n   E t h e r n e t - k a b e l . "  
 R B T _ U S B 	 = " U S B - a n s l u t n i n g "  
 H L P _ U S B 	 = " A n s l u t   % P R O D U C T % n   t i l l   e n   d a t o r   v i a   e n   U S B - k a b e l . "  
  
 [ W i f i A u t o C o n n e c t E r r o r ]  
 T I T L E 	 = " A u t o m a t i s k   W i - F i - a n s l u t n i n g   m i s s l y c k a d e s "  
 T I T L E _ W F D 	 = " T r � d l � s   a n s l u t n i n g   m i s s l y c k a d e s "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " A u t o m a t i s k   i n s t a l l a t i o n   a v   W i - F i   m i s s l y c k a d e s .   V � l j   e t t   a l t e r n a t i v   n e d a n   f � r   a t t   f o r t s � t t a   m e d   i n s t a l l a t i o n e n : \ r \ n 1 .   K l i c k a   p �   [ % B A C K % ]   f � r   a t t   f � r s � k a   i g e n .   \ r \ n 2 .   K l i c k a   p �   [ % N E X T % ]   f � r   a t t   a n s l u t a   t i l l   W i - F i   m e d   e n   a n n a n   m e t o d . "  
 T X T _ B o d y A P 	 = " I n s t � l l n i n g e n   h a r   m i s s l y c k a t s .   K l i c k a   p �   [ % B A C K % ]   o c h   f � r s � k   i g e n . "  
  
 [ I n f o r m a t i o n ]  
 T I T L E 	 = " V � l k o m m e n "  
 S U B _ T i t l e 	 = " T a c k   f � r   a t t   d u   h a r   v a l t   e n   E p s o n - % P R O D U C T % ! "  
 T X T _ C P 	 = " D u   k o m m e r   b l i   g u i d a d   g e n o m   i n s t a l l a t i o n s p r o c e s s e n   f � r   % P R O D U C T % n . "  
 T X T _ B P 	 = " P r o g r a m v a r a n   k o m m e r   a t t   i n s t a l l e r a s . "  
 T X T _ R e a d 	 = " N � r   % P R O D U C T % n   h a r   i n s t a l l e r a t s   k a n   d u   i n s t a l l e r a   y t t e r l i g a r e   p r o g r a m v a r a ,   t . e x .   u t s k r i f t s m � j l i g h e t e r   f � r   s u r f p l a t t a   e l l e r   s m a r t t e l e f o n . "  
  
 [ S S I D M a n u a l C o n n e c t ]  
 T I T L E 	 = " M a n u e l l   W i - F i - i n s t a l l a t i o n "  
 S U B _ T i t l e 	 = " "  
 I T M _ S S I D 	 = " N � t v e r k s n a m n   ( S S I D ) : "  
 I T M _ P W 	 = " L � s e n o r d : "  
 B T N _ S h o w P W 	 = " V i s a   l � s e n o r d "  
 I T M _ P W E r r o r 	 = " D e t   g i c k   i n t e   a t t   h � m t a "  
 I T M _ P W N o n e 	 = " O e t a b l e r a d "  
 L N K _ P u s h 	 = " I n s t a l l a t i o n   m e d   k n a p p t r y c k n i n g   f � r   W i - F i - n � t v e r k   ( W P S ) "  
  
 [ W i f i A u t o C o n n e c t ]  
 T I T L E 	 = " A u t o m a t i s k   W i - F i - i n s t a l l a t i o n "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D e t t a   u p p r � t t a r   a u t o m a t i s k t   e n   W i - F i - a n s l u t n i n g   t i l l   % P R O D U C T % n . "  
 C A U T I O N 	 = " I n t e r n e t a n s l u t n i n g e n   k o m m e r   a t t   i n a k t i v e r a s   t i l l f � l l i g t   m e d a n   e n   t r � d l � s   a n s l u t n i n g   u p p r � t t a s . \ r \ n S t � n g   a l l a   p r o g r a m   i n n a n   d u   s t a r t a r   i n s t a l l a t i o n e n . "  
 L N K _ S S I D 	 = " O m   d u   h e l l r e   v i l l   k o n f i g u r e r a   W i - F i - a n s l u t n i n g e n   m a n u e l l t   k l i c k a r   d u   h � r "  
 L N K _ W U S B 	 = " A u t o m a t i s k   i n s t a l l a t i o n   m e d   U S B - k a b e l "  
  
 [ E t h e r n e t C o n n e c t ]  
 T I T L E 	 = " E t h e r n e t - a n s l u t n i n g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " K o n t r o l l e r a   a t t   % P R O D U C T % n   � r   p �   o c h   a n s l u t   d e n   t i l l   r o u t e r n   m e d   e n   E t h e r n e t - k a b e l . "  
 C A U T I O N 	 = " K o n t r o l l e r a   a t t   d a t o r n   � r   a n s l u t e n   t i l l   n � t v e r k e t   ( a n t i n g e n   v i a   W i - F i   e l l e r   v i a   E t h e r n e t )   i n n a n   d u   f o r t s � t t e r . "  
  
 [ U S B W i r e d C o n n e c t ]  
 T I T L E 	 = " U S B - a n s l u t n i n g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " K o n t r o l l e r a   a t t   % P R O D U C T %   � r   p �   o c h   a n s l u t   d e n   t i l l   d a t o r n   v i a   e n   U S B - k a b e l . \ r \ n N � r   d a t o r n   h a r   h i t t a t   % P R O D U C T % n   v i s a s   n � s t a   s k � r m   a u t o m a t i s k t . "  
 C A U T I O N 	 = " "  
 C A U T I O N _ I F S 	 = " S t � l l   i n   o m k o p p l a r e n s   a n s l u t n i n g s l � g e   p �   p r o d u k t e n   t i l l   U S B ,   o c h   a n s l u t   s e d a n   U S B - k a b e l n . "  
 C B X _ L a t e r 	 = " A n s l u t   % P R O D U C T % n   v i d   e t t   s e n a r e   t i l l f � l l e "  
  
 [ W i f i A u t o C o n n e c t W i t h U S B ]  
 T I T L E 	 = " A u t o m a t i s k   W i - F i - i n s t a l l a t i o n   ( t i l l f � l l i g   a n v � n d n i n g   a v   e n   U S B - k a b e l ) "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " K o n t r o l l e r a   a t t   % P R O D U C T % n   � r   p �   o c h   a n s l u t   d e n   t i l l   d a t o r n   v i a   e n   U S B - k a b e l   ( d u   b e h � v e r   b a r a   t i l l f � l l i g t   a n s l u t a   U S B - k a b e l n   u n d e r   W i - F i - i n s t a l l a t i o n e n ) .   \ r \ n N � r   d a t o r n   h i t t a r   % P R O D U C T % n   v i s a s   n � s t a   s k � r m   a u t o m a t i s k t . "  
 C A U T I O N 	 = " K o p p l a   i n t e   u r   U S B - k a b e l n   f � r r � n   d u   o m b e d s   g � r a   d e t . "  
 L N K _ P U S H 	 = " I n s t a l l a t i o n   m e d   k n a p p t r y c k n i n g   f � r   W i - F i - n � t v e r k   ( W P S ) "  
  
 [ W i f i D i r e c t C o n n e c t ]  
 T I T L E 	 = " A n s l u t n i n g   m e d   W i - F i   D i r e c t "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D e t   h � r   u p p r � t t a r   e n   d i r e k t   W i - F i - a n s l u t n i n g   m e l l a n   d a t o r n   o c h   % P R O D U C T % n . \ r \ n S e   b r u k s a n v i s n i n g e n   f � r   m e r   i n f o r m a t i o n   o m   W i - F i   D i r e c t . "  
 C A U T I O N 	 = " V i   r e k o m m e n d e r a r   i n t e   d e n   h � r   a n s l u t n i n g s m e t o d e n   o m   d u   h a r   e n   W i - F i - r o u t e r . "  
  
 [ D i r e c t W i f i C o n n e c t ]  
 T I T L E 	 = " S t � l l   i n   d i r e k t   W i - F i - a n s l u t n i n g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D e t t a   s k a p a r   e n   d i r e k t   W i - F i - a n s l u t n i n g   m e l l a n   d e n   h � r   d a t o r n   o c h   % P R O D U C T % . \ r \ n S e   h a n d b o k e n   f � r   y t t e r l i g a r e   i n f o r m a t i o n   o m   d i r e k t   W i - F i - a n s l u t n i n g . "  
 C A U T I O N 	 = " V i   r e k o m m e n d e r a r   i n t e   d e n   h � r   a n s l u t n i n g s m e t o d e n   o m   d u   h a r   e n   W i - F i - r o u t e r . "  
  
 [ W F D M a n u a l ]  
 T I T L E 	 = " I n s t � l l n i n g   f � r   t r � d l � s   a n s l u t n i n g s h a n d b o k "  
 S U B _ T i t l e 	 = " "  
  
 [ P u s h B u t t o n C o n n e c t ]  
 T I T L E 	 = " I n s t a l l a t i o n   m e d   k n a p p t r y c k n i n g   f � r   W i - F i - n � t v e r k   ( W P S ) "  
 S U B _ T i t l e 	 = " "  
 L N K _ A P m o d e 	 = " K l i c k a   h � r   o m   d i n   t r � d l � s a   r o u t e r   i n t e   s t � d e r   W P S - t r y c k k n a p p s f u n k t i o n e n "  
  
 [ A P m o d e M a n u a l S e t t i n g ]  
 T I T L E                 = " I n s t � l l n i n g   f � r   t r � d l � s   a n s l u t n i n g s h a n d b o k "  
  
 [ I P M a n u a l C o n n e c t ]  
 T I T L E 	 = " I n s t � l l n i n g   a v   n � t v e r k s p o r t "  
 S U B _ T i t l e 	 = " "  
 T X T _ S e t t i n g 	 = " S t � l l e r   i n   a n s l u t n i n g . . .   v � n t a . "  
  
 [ I n s t a l l N e t w o r k ]  
 T I T L E 	 = " I n s t a l l e r a r   n � t v e r k s v e r k t y g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y _ D L 	 = " H � m t a r   . . .   % s "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   . . .   % s "  
  
 [ N e t w o r k C o n n e c t e d ]  
 T I T L E 	 = " I n s t a l l a t i o n e n   � r   k l a r "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " P r o g r a m v a r u -   o c h   n � t v e r k s i n s t a l l a t i o n e n   h a r   s l u t f � r t s . "  
 S P I N F O 	 = " K o p p l a   u r   U S B - k a b e l n   o m   d u   h a r   a n v � n t   d e n   t i l l   n � t v e r k s i n s t a l l a t i o n e n . "  
 I T M _ P r i n t e r 	 = " S k r i v a r d r i v r u t i n "  
 I T M _ P o r t 	 = " P o r t n a m n "  
 I T M _ I P A d d r e s s 	 = " I P - a d r e s s "  
 I T M _ M a c A d d r e s s 	 = " M A C - a d r e s s "  
  
 [ L o c a l C o n n e c t e d ]  
 T I T L E 	 = " I n s t a l l a t i o n e n   � r   k l a r "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " P r o g r a m v a r u i n s t a l l a t i o n e n   v i a   U S B   h a r   s l u t f � r t s . "  
 I T M _ P r i n t e r 	 = " S k r i v a r d r i v r u t i n "  
 I T M _ P o r t 	 = " P o r t n a m n "  
  
 [ W a i t I n i t i a l C h a r g e ]  
 T I T L E               = " S t a r t a r . . . "  
 T X T _ B o d y   = " B l � c k s y s t e m e t   s t a r t a r . . . v a r   g o d   v � n t a . "  
  
 [ T e s t P r i n t ]  
 T I T L E 	 = " S k r i v   u t   t e s t s i d a "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " K l i c k a   p �   [ % P R I N T % ]   f � r   a t t   k o n t r o l l e r a   a t t   i n s t a l l a t i o n e n   a v   p r o g r a m v a r a   o c h   k o n f i g u r a t i o n e n   a v   % P R O D U C T %   h a r   s l u t f � r t s . "  
 L N K _ U t i l l i t y 	 = " K l i c k a   h � r   o m   u t s k r i f t s k v a l i t e t e n   � r   d � l i g . "  
 B T N _ P r i n t 	 = " S k r i v   u t   t e s t s i d a "  
  
 [ I n v i t a t i o n ]  
 T I T L E 	 = " P r o d u k t r e g i s t r e r i n g   o n l i n e "  
 S U B _ T i t l e _ P R O D U C T 	 = " P r o d u k t n a m n "  
 S U B _ T i t l e _ S E R I A L 	 = " S e r i e n u m m e r "  
 R B T _ I n s t a l l 	 = " I n s t a l l e r a "  
 R B T _ D i s a g r e e 	 = " I n s t a l l e r a   i n t e "  
 R B T _ L a t e r 	 = " P � m i n n   m i g   s e n a r e "  
 T X T _ L o a d i n g 	 = " L a d d a r . . . "  
 T X T _ B o d y _ D L 	 = " H � m t a r   . . .   % s "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   . . .   % s "  
 T X T _ R e g i o n 	 = " V � l j   d i t t   l a n d / r e g i o n . "  
 T X T _ N W _ E r r o r 	 = " K a n   i n t e   a n s l u t a   t i l l   i n t e r n e t .   K o n t r o l l e r a   d i n   a n s l u t n i n g   o c h   f � r s � k   i g e n . "  
  
 [ W a r r a n t y ]  
 T I T L E 	 	 = " I s s u e   r e q u e s t i n g   t h e   w a r r a n t y   c a r d   a n d   o n l i n e   p r o d u c t   r e g i s t r a t i o n "  
 S U B _ T i t l e 	 = " "  
 I T M _ P R O D U C T 	 = " P r o d u k t n a m n "  
 I T M _ S E R I A L 	 = " S e r i e n u m m e r "  
 I T M _ E R E G 	 	 = " P r o d u k t r e g i s t r e r i n g   o n l i n e "  
 T X T _ E R E G _ M E S S A G E 	 = " T h i s   p r o d u c t   c a n   p e r f o r m   o n l i n e   u s e r   r e g i s t r a t i o n .   \ r \ n W h e n   y o u   r e g i s t e r ,   y o u   r e c e i v e   f r o m   a   d e d i c a t e d   s i t e   o r   e - m a i l ,   a n d   r e l a t e d   i n f o r m a t i o n ,   s u c h   a s   s o f t w a r e   u p d a t e s   a n d   d r i v e r s   i n f o r m a t i o n   o f   t h e   p r o d u c t . "  
 I T M _ W A R R A N T Y 	 = " I s s u e   r e q u e s t i n g   t h e   w a r r a n t y   c a r d "  
 T X T W A R R A N T Y _ M E S S A G E 	 = " Y o u   c a n   r e q u e s t   b y   m a i l   o r   W e b . "  
 T X T _ B U T T O N _ M E S S A G E 	 = " I f   y o u   w a n t   t o   i s s u e   c l a i m s   o f   w a r r a n t y   c a r d   a n d   p r o d u c t   r e g i s t r a t i o n ,   p l e a s e   c l i c k   [ W a r r a n t y   c a r d   r e q u e s t   /   O n l i n e   r e g i s t r a t i o n ] . \ r \ n I f   y o u   o n l y   w a n t   t o   i s s u e   c l a i m s   w a r r a n t y   c a r d ,   p l e a s e   c l i c k   [ W a r r a n t y   c a r d   r e q u e s t ] . "  
 B T N _ E R E G 	 	 = " W a r r a n t y   c a r d   r e q u e s t   /   O n l i n e   r e g i s t r a t i o n "  
 B T N _ W A R R A N T Y 	 = " W a r r a n t y   c a r d   r e q u e s t "  
 T X T _ M E S S A G E _ M U L T = " Y o u   c a n   r e g i s t e r   t h e   p r o d u c t   s e l e c t i o n   i s   n o t   i n   t h e   s e r i a l   n u m b e r   f i e l d . "  
 T X T _ M E S S A G E _ O N E 	 = " Y o u   c a n   r e g i s t e r   t h e   p r o d u c t   d i f f e r e n t   f r o m   w h a t   y o u   s e e   o n   y o u r   s e r i a l   n u m b e r   f i e l d . "  
 T X T _ N W _ E R R O R 	 = " Y o u   c a n   n o t   c o n n e c t   t o   t h e   I n t e r n e t .   O n   t h e   c h e c k ,   p l e a s e   t r y   a g a i n   t h e   c o n n e c t i o n   s t a t u s   t o   t h e   I n t e r n e t . \ r \ n I f   y o u   c a n   n o t   c o n n e c t   t o   t h e   I n t e r n e t ,   p l e a s e   a p p l y   b y   w a r r a n t y   c a r d   i s s u e d   r e q u e s t   f o r m   t h a t   i s   i n c l u d e d   i n   t h e   p r o d u c t . "  
  
  
 [ F i n i s h ]  
 T I T L E 	 = " E x t r a p r o g r a m "  
 T I T L E _ N o S W 	 = " I n s t a l l a t i o n e n   � r   k l a r "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " P �   f � l j a n d e   s k � r m   k a n   d u   v � l j a   a t t   i n s t a l l e r a   � v r i g   p r o g r a m v a r a   s o m . "  
 T X T _ R e a d 	 = " -   U t s k r i f t s m � j l i g h e t   f r � n   s m a r t t e l e f o n   o c h   s u r f p l a t t a \ r \ n -   V i k t i g a   u p p d a t e r i n g a r   f � r   % P R O D U C T % n   \ r \ n -   U t s k r i f t s -   o c h   s k a n n i n g s a p p a r   f r � n   E p s o n "  
  
 [ S y s t e m E r r o r ]  
 T I T L E 	 = " S y s t e m f e l "  
 E R R _ A d m i n 	 = " D u   m � s t e   v a r a   i n l o g g a d   s o m   a d m i n i s t r a t � r   f � r   a t t   k u n n a   i n s t a l l e r a   p r o g r a m v a r a n . "  
 E R R _ O S 	 = " D i t t   o p e r a t i v s y s t e m   h a r   i n t e   s t � d   f � r   p r o g r a m v a r a n . "  
 E R R _ H D D 	 = " D e t   f i n n s   i n t e   t i l l r � c k l i g t   m e d   l e d i g t   u t r y m m e . \ r \ n V � l j   a t t   i n s t a l l e r a   f � r r e   o b j e k t   e l l e r   f r i g � r   m e r   u t r y m m e   o c h   i n s t a l l e r a   p r o g r a m v a r a n   i g e n . "  
  
 [ N W S e t t i n g E r r o r ]  
 T I T L E 	 = " N � t v e r k s k o n f i g u r a t i o n e n   a v b r � t s "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
 T X T _ R e s t a r t 	 = " P r o d u k t n a m n e t   s o m   d u   h a r   v a l t   k a n   v a r a   f e l . "  
  
 [ T i m e O u t E r r o r ]  
 T I T L E 	 = " % P R O D U C T % n   k � n n s   i n t e   i g e n "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
 T X T _ R e s t a r t 	 = " P r o d u k t n a m n e t   s o m   d u   h a r   v a l t   k a n   v a r a   f e l . "  
  
 [ A b n o m a l E r r o r ]  
 T I T L E 	 = " F e l   v i d   a n s l u t n i n g   t i l l   n � t v e r k "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
  
 [ W a i t C o n n e c t ]  
 T I T L E 	 = " N � t v e r k s k o n f i g u r a t i o n "  
 S U B _ T i t l e 	 = " H � m t a r   E p s o n N e t   S e t u p "  
 T X T _ B o d y 	 = " V � n t a   . . . "  
  
 [ W a i t S o f t w a r e ]  
 T I T L E 	 = " I n s t a l l e r a   t i l l � m p n i n g s p r o g r a m "  
 S U B _ T i t l e 	 = " A n s l u t e r   t i l l   E p s o n   S o f t w a r e   U p d a t e r "  
 T X T _ B o d y 	 = " V � n t a   . . . "  
  
 [ N e t w o r k E r r o r ]  
 T I T L E 	 = " F e l   v i d   a n s l u t n i n g   t i l l   n � t v e r k "  
 S U B _ T i t l e 	 = " N � t v e r k e t s   g r � n s s n i t t   � r   i n t e   t i l l g � n g l i g t . "  
  
 [ W e b D o w n l o a d E r r o r ]  
 T I T L E 	 = " F e l   v i d   h � m t n i n g   a v   f i l "  
 E R R _ F a i l e d 	 = " D e t   g i c k   i n t e   a t t   a n s l u t a   t i l l   I n t e r n e t .   K o n t r o l l e r a   d i n   I n t e r n e t a n s l u t n i n g . "  
 E R R _ C o m m 	 = " D e t   g i c k   i n t e   a t t   a n s l u t a   t i l l   I n t e r n e t .   K o n t r o l l e r a   d i n   I n t e r n e t a n s l u t n i n g . "  
  
 [ S o f t w a r e N a m e ]  
 P r i n t e r D r i v e r x 6 4 	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 6 4 _ L P 	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 _ L P 	 = " S k r i v a r d r i v r u t i n "  
 S c a n n e r D r i v e r 	 = " S k a n n e r d r i v r u t i n "  
 I S I S D r i v e r 	 = " E M C   I S I S   D r i v e r "  
 E p s o n N e t P r i n t E 	 = " E p s o n N e t   P r i n t "  
 E p s o n N e t P r i n t J 	 = " E p s o n N e t   P r i n t "  
 E p s o n S c a n O C R C o m p o n e n t 	 = " E p s o n   S c a n   O C R   C o m p o n e n t "  
 E p s o n S c a n P D F E x t e n s i o n s 	 = " E p s o n   S c a n   P D F   E x t e n s i o n s "  
 E v e n t M a n a g e r 	 = " E v e n t   M a n a g e r "  
 D o c u m e n t C a p t u r e 	 = " D o c u m e n t   C a p t u r e   P r o "  
 M y E P S O N P o r t a l 	 = " M y E P S O N   P o r t a l "  
 D o w n l o a d N a v i g a t o r 	 = " S o f t w a r e   U p d a t e r "  
 E p s o n N e t S e t u p 	 = " E p s o n N e t   S e t u p "  
 E p s o n N e t C o n f i g 	 = " E p s o n N e t   C o n f i g "  
 M a n u a l P a c k a g e 	 = " E p s o n   M a n u a l   P a c k a g e "  
 E p s o n C o n n e c t S h o r t c u t 	 = " E p s o n   C o n n e c t   S i t e "  
 F a x U t i l i t y 	 = " F a x   U t i l i t y "  
 F a x U t i l i t y W 	 = " F a x   U t i l i t y "  
 P I F I n s t a l l e r 	 = " P R I N T   I m a g e   F r a m e r "  
 B u s i n e s s C a r d F i l i n g E n t r y 	 = " B u s i n e s s   C a r d   F i l i n g   E n t r y "  
 